module Mux4(in0,in1,in2,in3,out,src);
input [31:0] in0, in1, in2, in3;
input [1:0] src;
output reg [31:0] out;

always @(src or in0 or in1 or in2 or in3) begin
    case(src)
    2'b00: out <= in0;
    2'b01: out <= in1;
    2'b10: out <= in2;
    2'b11: out <= in3;
    endcase
end
endmodule